`include "hazard_unit_if.vh"

module hazard_unit(hazard_unit_if.hu huif);
endmodule
