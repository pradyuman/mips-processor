`include "forwarding_unit_if.vh"

module forwarding_unit(forwarding_unit_if.fu fuif);
endmodule
